--BIBLIOTECAS USADAS PARA REALIZAÇÃO DO PROGRAMA
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity teste0 is
	port
	(
	   -- ENTRADAS FISICAS!
		-- Obs:Não existe necessidade de modificar nada aqui!!!
		
		--DE0Nano
		-- Input ports 
		CLOCK_50 : in std_logic; -- Oscilador
		KEY : in std_logic_vector( 1 downto 0); --Botões que ficam na placa DE0-nano
		
		--output ports
		LED : out std_logic_vector(2 downto 0); --LEDS que ficam na placa DEO-nano

		--Expansion Header UFPE/DES kit
		-- input ports
		ehkey : in std_logic_vector(4 downto 0);-- bits 0-7=>chaves; bits 8 e 9 => pushbutton
		
		-- output ports
		dig7seg : out std_logic_vector(1 downto 0); -- Seletor do display
		d7seg : out std_logic_vector(8 downto 0) -- Indicator de 7seg selecionado por dig7seg
		
	);
end teste0;


architecture behaviorOfTest of teste0 is
--Colocar aqui todas os sinais que deseja utilizar("equivalentes a variaveis auxiliares")
signal vtest: std_logic_vector(4 downto 0);
begin

process(clock_50) -- Divisor do sinal de clock da placa(50Mhz)
variable count: integer range 0 to 50000000;
begin
	if rising_edge(clock_50) then
		count:=count+1;
		if count=(20*2500000) then
			count:=0;
			if unsigned(vtest)>=9 then
				vtest<=(others=>'0');
			else
				vtest<=std_logic_vector(unsigned(vtest)+1);
			end if;
		end if;
	end if;
end process;


LED(4 downto 0)<=vtest;
 
end behaviorOfTest;
